`timescale 1ps/1ps